/////////////////////////////////////////////////////////////////////
//
//
//Author : Elsie Rezinold Yedida
//
//
//
/////////////////////////////////////////////////////////////////////







module dm (
    clk,
    rst_n,
    i_byte_rd,
    i_2byte_rd,
    i_4byte_rd,
    i_mem_rd,
    i_se_mem_rd,
    i_address,
    o_rd_data,
    i_byte_wr,
    i_2byte_wr,
    i_4byte_wr,
    i_mem_wr,
    i_wr_data
);


input [0:0] clk;
input rst_n;
input [0:0] i_byte_rd;
input [0:0] i_2byte_rd;
input [0:0] i_4byte_rd;
input [0:0] i_mem_rd;
input [0:0] i_se_mem_rd;
input [31:0] i_address;
output [31:0] o_rd_data;
input [0:0] i_byte_wr;
input [0:0] i_2byte_wr;
input [0:0] i_4byte_wr;
input [0:0] i_mem_wr;
input [31:0] i_wr_data;

reg [31:0] w_rd_data;
reg [15:0] w_rd_data_2byte;
reg [7:0] w_rd_data_byte;
reg [31:0] mem [0:1024-1];



always @(posedge clk, negedge rst_n) begin
    if (rst_n == 0) begin
        mem[0] <= 0;
        mem[1] <= 0;
        mem[2] <= 0;
        mem[3] <= 0;
        mem[4] <= 0;
        mem[5] <= 0;
        mem[6] <= 0;
        mem[7] <= 0;
        mem[8] <= 0;
        mem[9] <= 0;
        mem[10] <= 0;
        mem[11] <= 0;
        mem[12] <= 0;
        mem[13] <= 0;
        mem[14] <= 0;
        mem[15] <= 0;
        mem[16] <= 0;
        mem[17] <= 0;
        mem[18] <= 0;
        mem[19] <= 0;
        mem[20] <= 0;
        mem[21] <= 0;
        mem[22] <= 0;
        mem[23] <= 0;
        mem[24] <= 0;
        mem[25] <= 0;
        mem[26] <= 0;
        mem[27] <= 0;
        mem[28] <= 0;
        mem[29] <= 0;
        mem[30] <= 0;
        mem[31] <= 0;
        mem[32] <= 0;
        mem[33] <= 0;
        mem[34] <= 0;
        mem[35] <= 0;
        mem[36] <= 0;
        mem[37] <= 0;
        mem[38] <= 0;
        mem[39] <= 0;
        mem[40] <= 0;
        mem[41] <= 0;
        mem[42] <= 0;
        mem[43] <= 0;
        mem[44] <= 0;
        mem[45] <= 0;
        mem[46] <= 0;
        mem[47] <= 0;
        mem[48] <= 0;
        mem[49] <= 0;
        mem[50] <= 0;
        mem[51] <= 0;
        mem[52] <= 0;
        mem[53] <= 0;
        mem[54] <= 0;
        mem[55] <= 0;
        mem[56] <= 0;
        mem[57] <= 0;
        mem[58] <= 0;
        mem[59] <= 0;
        mem[60] <= 0;
        mem[61] <= 0;
        mem[62] <= 0;
        mem[63] <= 0;
        mem[64] <= 0;
        mem[65] <= 0;
        mem[66] <= 0;
        mem[67] <= 0;
        mem[68] <= 0;
        mem[69] <= 0;
        mem[70] <= 0;
        mem[71] <= 0;
        mem[72] <= 0;
        mem[73] <= 0;
        mem[74] <= 0;
        mem[75] <= 0;
        mem[76] <= 0;
        mem[77] <= 0;
        mem[78] <= 0;
        mem[79] <= 0;
        mem[80] <= 0;
        mem[81] <= 0;
        mem[82] <= 0;
        mem[83] <= 0;
        mem[84] <= 0;
        mem[85] <= 0;
        mem[86] <= 0;
        mem[87] <= 0;
        mem[88] <= 0;
        mem[89] <= 0;
        mem[90] <= 0;
        mem[91] <= 0;
        mem[92] <= 0;
        mem[93] <= 0;
        mem[94] <= 0;
        mem[95] <= 0;
        mem[96] <= 0;
        mem[97] <= 0;
        mem[98] <= 0;
        mem[99] <= 0;
        mem[100] <= 0;
        mem[101] <= 0;
        mem[102] <= 0;
        mem[103] <= 0;
        mem[104] <= 0;
        mem[105] <= 0;
        mem[106] <= 0;
        mem[107] <= 0;
        mem[108] <= 0;
        mem[109] <= 0;
        mem[110] <= 0;
        mem[111] <= 0;
        mem[112] <= 0;
        mem[113] <= 0;
        mem[114] <= 0;
        mem[115] <= 0;
        mem[116] <= 0;
        mem[117] <= 0;
        mem[118] <= 0;
        mem[119] <= 0;
        mem[120] <= 0;
        mem[121] <= 0;
        mem[122] <= 0;
        mem[123] <= 0;
        mem[124] <= 0;
        mem[125] <= 0;
        mem[126] <= 0;
        mem[127] <= 0;
        mem[128] <= 0;
        mem[129] <= 0;
        mem[130] <= 0;
        mem[131] <= 0;
        mem[132] <= 0;
        mem[133] <= 0;
        mem[134] <= 0;
        mem[135] <= 0;
        mem[136] <= 0;
        mem[137] <= 0;
        mem[138] <= 0;
        mem[139] <= 0;
        mem[140] <= 0;
        mem[141] <= 0;
        mem[142] <= 0;
        mem[143] <= 0;
        mem[144] <= 0;
        mem[145] <= 0;
        mem[146] <= 0;
        mem[147] <= 0;
        mem[148] <= 0;
        mem[149] <= 0;
        mem[150] <= 0;
        mem[151] <= 0;
        mem[152] <= 0;
        mem[153] <= 0;
        mem[154] <= 0;
        mem[155] <= 0;
        mem[156] <= 0;
        mem[157] <= 0;
        mem[158] <= 0;
        mem[159] <= 0;
        mem[160] <= 0;
        mem[161] <= 0;
        mem[162] <= 0;
        mem[163] <= 0;
        mem[164] <= 0;
        mem[165] <= 0;
        mem[166] <= 0;
        mem[167] <= 0;
        mem[168] <= 0;
        mem[169] <= 0;
        mem[170] <= 0;
        mem[171] <= 0;
        mem[172] <= 0;
        mem[173] <= 0;
        mem[174] <= 0;
        mem[175] <= 0;
        mem[176] <= 0;
        mem[177] <= 0;
        mem[178] <= 0;
        mem[179] <= 0;
        mem[180] <= 0;
        mem[181] <= 0;
        mem[182] <= 0;
        mem[183] <= 0;
        mem[184] <= 0;
        mem[185] <= 0;
        mem[186] <= 0;
        mem[187] <= 0;
        mem[188] <= 0;
        mem[189] <= 0;
        mem[190] <= 0;
        mem[191] <= 0;
        mem[192] <= 0;
        mem[193] <= 0;
        mem[194] <= 0;
        mem[195] <= 0;
        mem[196] <= 0;
        mem[197] <= 0;
        mem[198] <= 0;
        mem[199] <= 0;
        mem[200] <= 0;
        mem[201] <= 0;
        mem[202] <= 0;
        mem[203] <= 0;
        mem[204] <= 0;
        mem[205] <= 0;
        mem[206] <= 0;
        mem[207] <= 0;
        mem[208] <= 0;
        mem[209] <= 0;
        mem[210] <= 0;
        mem[211] <= 0;
        mem[212] <= 0;
        mem[213] <= 0;
        mem[214] <= 0;
        mem[215] <= 0;
        mem[216] <= 0;
        mem[217] <= 0;
        mem[218] <= 0;
        mem[219] <= 0;
        mem[220] <= 0;
        mem[221] <= 0;
        mem[222] <= 0;
        mem[223] <= 0;
        mem[224] <= 0;
        mem[225] <= 0;
        mem[226] <= 0;
        mem[227] <= 0;
        mem[228] <= 0;
        mem[229] <= 0;
        mem[230] <= 0;
        mem[231] <= 0;
        mem[232] <= 0;
        mem[233] <= 0;
        mem[234] <= 0;
        mem[235] <= 0;
        mem[236] <= 0;
        mem[237] <= 0;
        mem[238] <= 0;
        mem[239] <= 0;
        mem[240] <= 0;
        mem[241] <= 0;
        mem[242] <= 0;
        mem[243] <= 0;
        mem[244] <= 0;
        mem[245] <= 0;
        mem[246] <= 0;
        mem[247] <= 0;
        mem[248] <= 0;
        mem[249] <= 0;
        mem[250] <= 0;
        mem[251] <= 0;
        mem[252] <= 0;
        mem[253] <= 0;
        mem[254] <= 0;
        mem[255] <= 0;
        mem[256] <= 0;
        mem[257] <= 0;
        mem[258] <= 0;
        mem[259] <= 0;
        mem[260] <= 0;
        mem[261] <= 0;
        mem[262] <= 0;
        mem[263] <= 0;
        mem[264] <= 0;
        mem[265] <= 0;
        mem[266] <= 0;
        mem[267] <= 0;
        mem[268] <= 0;
        mem[269] <= 0;
        mem[270] <= 0;
        mem[271] <= 0;
        mem[272] <= 0;
        mem[273] <= 0;
        mem[274] <= 0;
        mem[275] <= 0;
        mem[276] <= 0;
        mem[277] <= 0;
        mem[278] <= 0;
        mem[279] <= 0;
        mem[280] <= 0;
        mem[281] <= 0;
        mem[282] <= 0;
        mem[283] <= 0;
        mem[284] <= 0;
        mem[285] <= 0;
        mem[286] <= 0;
        mem[287] <= 0;
        mem[288] <= 0;
        mem[289] <= 0;
        mem[290] <= 0;
        mem[291] <= 0;
        mem[292] <= 0;
        mem[293] <= 0;
        mem[294] <= 0;
        mem[295] <= 0;
        mem[296] <= 0;
        mem[297] <= 0;
        mem[298] <= 0;
        mem[299] <= 0;
        mem[300] <= 0;
        mem[301] <= 0;
        mem[302] <= 0;
        mem[303] <= 0;
        mem[304] <= 0;
        mem[305] <= 0;
        mem[306] <= 0;
        mem[307] <= 0;
        mem[308] <= 0;
        mem[309] <= 0;
        mem[310] <= 0;
        mem[311] <= 0;
        mem[312] <= 0;
        mem[313] <= 0;
        mem[314] <= 0;
        mem[315] <= 0;
        mem[316] <= 0;
        mem[317] <= 0;
        mem[318] <= 0;
        mem[319] <= 0;
        mem[320] <= 0;
        mem[321] <= 0;
        mem[322] <= 0;
        mem[323] <= 0;
        mem[324] <= 0;
        mem[325] <= 0;
        mem[326] <= 0;
        mem[327] <= 0;
        mem[328] <= 0;
        mem[329] <= 0;
        mem[330] <= 0;
        mem[331] <= 0;
        mem[332] <= 0;
        mem[333] <= 0;
        mem[334] <= 0;
        mem[335] <= 0;
        mem[336] <= 0;
        mem[337] <= 0;
        mem[338] <= 0;
        mem[339] <= 0;
        mem[340] <= 0;
        mem[341] <= 0;
        mem[342] <= 0;
        mem[343] <= 0;
        mem[344] <= 0;
        mem[345] <= 0;
        mem[346] <= 0;
        mem[347] <= 0;
        mem[348] <= 0;
        mem[349] <= 0;
        mem[350] <= 0;
        mem[351] <= 0;
        mem[352] <= 0;
        mem[353] <= 0;
        mem[354] <= 0;
        mem[355] <= 0;
        mem[356] <= 0;
        mem[357] <= 0;
        mem[358] <= 0;
        mem[359] <= 0;
        mem[360] <= 0;
        mem[361] <= 0;
        mem[362] <= 0;
        mem[363] <= 0;
        mem[364] <= 0;
        mem[365] <= 0;
        mem[366] <= 0;
        mem[367] <= 0;
        mem[368] <= 0;
        mem[369] <= 0;
        mem[370] <= 0;
        mem[371] <= 0;
        mem[372] <= 0;
        mem[373] <= 0;
        mem[374] <= 0;
        mem[375] <= 0;
        mem[376] <= 0;
        mem[377] <= 0;
        mem[378] <= 0;
        mem[379] <= 0;
        mem[380] <= 0;
        mem[381] <= 0;
        mem[382] <= 0;
        mem[383] <= 0;
        mem[384] <= 0;
        mem[385] <= 0;
        mem[386] <= 0;
        mem[387] <= 0;
        mem[388] <= 0;
        mem[389] <= 0;
        mem[390] <= 0;
        mem[391] <= 0;
        mem[392] <= 0;
        mem[393] <= 0;
        mem[394] <= 0;
        mem[395] <= 0;
        mem[396] <= 0;
        mem[397] <= 0;
        mem[398] <= 0;
        mem[399] <= 0;
        mem[400] <= 0;
        mem[401] <= 0;
        mem[402] <= 0;
        mem[403] <= 0;
        mem[404] <= 0;
        mem[405] <= 0;
        mem[406] <= 0;
        mem[407] <= 0;
        mem[408] <= 0;
        mem[409] <= 0;
        mem[410] <= 0;
        mem[411] <= 0;
        mem[412] <= 0;
        mem[413] <= 0;
        mem[414] <= 0;
        mem[415] <= 0;
        mem[416] <= 0;
        mem[417] <= 0;
        mem[418] <= 0;
        mem[419] <= 0;
        mem[420] <= 0;
        mem[421] <= 0;
        mem[422] <= 0;
        mem[423] <= 0;
        mem[424] <= 0;
        mem[425] <= 0;
        mem[426] <= 0;
        mem[427] <= 0;
        mem[428] <= 0;
        mem[429] <= 0;
        mem[430] <= 0;
        mem[431] <= 0;
        mem[432] <= 0;
        mem[433] <= 0;
        mem[434] <= 0;
        mem[435] <= 0;
        mem[436] <= 0;
        mem[437] <= 0;
        mem[438] <= 0;
        mem[439] <= 0;
        mem[440] <= 0;
        mem[441] <= 0;
        mem[442] <= 0;
        mem[443] <= 0;
        mem[444] <= 0;
        mem[445] <= 0;
        mem[446] <= 0;
        mem[447] <= 0;
        mem[448] <= 0;
        mem[449] <= 0;
        mem[450] <= 0;
        mem[451] <= 0;
        mem[452] <= 0;
        mem[453] <= 0;
        mem[454] <= 0;
        mem[455] <= 0;
        mem[456] <= 0;
        mem[457] <= 0;
        mem[458] <= 0;
        mem[459] <= 0;
        mem[460] <= 0;
        mem[461] <= 0;
        mem[462] <= 0;
        mem[463] <= 0;
        mem[464] <= 0;
        mem[465] <= 0;
        mem[466] <= 0;
        mem[467] <= 0;
        mem[468] <= 0;
        mem[469] <= 0;
        mem[470] <= 0;
        mem[471] <= 0;
        mem[472] <= 0;
        mem[473] <= 0;
        mem[474] <= 0;
        mem[475] <= 0;
        mem[476] <= 0;
        mem[477] <= 0;
        mem[478] <= 0;
        mem[479] <= 0;
        mem[480] <= 0;
        mem[481] <= 0;
        mem[482] <= 0;
        mem[483] <= 0;
        mem[484] <= 0;
        mem[485] <= 0;
        mem[486] <= 0;
        mem[487] <= 0;
        mem[488] <= 0;
        mem[489] <= 0;
        mem[490] <= 0;
        mem[491] <= 0;
        mem[492] <= 0;
        mem[493] <= 0;
        mem[494] <= 0;
        mem[495] <= 0;
        mem[496] <= 0;
        mem[497] <= 0;
        mem[498] <= 0;
        mem[499] <= 0;
        mem[500] <= 0;
        mem[501] <= 0;
        mem[502] <= 0;
        mem[503] <= 0;
        mem[504] <= 0;
        mem[505] <= 0;
        mem[506] <= 0;
        mem[507] <= 0;
        mem[508] <= 0;
        mem[509] <= 0;
        mem[510] <= 0;
        mem[511] <= 0;
        mem[512] <= 0;
        mem[513] <= 0;
        mem[514] <= 0;
        mem[515] <= 0;
        mem[516] <= 0;
        mem[517] <= 0;
        mem[518] <= 0;
        mem[519] <= 0;
        mem[520] <= 0;
        mem[521] <= 0;
        mem[522] <= 0;
        mem[523] <= 0;
        mem[524] <= 0;
        mem[525] <= 0;
        mem[526] <= 0;
        mem[527] <= 0;
        mem[528] <= 0;
        mem[529] <= 0;
        mem[530] <= 0;
        mem[531] <= 0;
        mem[532] <= 0;
        mem[533] <= 0;
        mem[534] <= 0;
        mem[535] <= 0;
        mem[536] <= 0;
        mem[537] <= 0;
        mem[538] <= 0;
        mem[539] <= 0;
        mem[540] <= 0;
        mem[541] <= 0;
        mem[542] <= 0;
        mem[543] <= 0;
        mem[544] <= 0;
        mem[545] <= 0;
        mem[546] <= 0;
        mem[547] <= 0;
        mem[548] <= 0;
        mem[549] <= 0;
        mem[550] <= 0;
        mem[551] <= 0;
        mem[552] <= 0;
        mem[553] <= 0;
        mem[554] <= 0;
        mem[555] <= 0;
        mem[556] <= 0;
        mem[557] <= 0;
        mem[558] <= 0;
        mem[559] <= 0;
        mem[560] <= 0;
        mem[561] <= 0;
        mem[562] <= 0;
        mem[563] <= 0;
        mem[564] <= 0;
        mem[565] <= 0;
        mem[566] <= 0;
        mem[567] <= 0;
        mem[568] <= 0;
        mem[569] <= 0;
        mem[570] <= 0;
        mem[571] <= 0;
        mem[572] <= 0;
        mem[573] <= 0;
        mem[574] <= 0;
        mem[575] <= 0;
        mem[576] <= 0;
        mem[577] <= 0;
        mem[578] <= 0;
        mem[579] <= 0;
        mem[580] <= 0;
        mem[581] <= 0;
        mem[582] <= 0;
        mem[583] <= 0;
        mem[584] <= 0;
        mem[585] <= 0;
        mem[586] <= 0;
        mem[587] <= 0;
        mem[588] <= 0;
        mem[589] <= 0;
        mem[590] <= 0;
        mem[591] <= 0;
        mem[592] <= 0;
        mem[593] <= 0;
        mem[594] <= 0;
        mem[595] <= 0;
        mem[596] <= 0;
        mem[597] <= 0;
        mem[598] <= 0;
        mem[599] <= 0;
        mem[600] <= 0;
        mem[601] <= 0;
        mem[602] <= 0;
        mem[603] <= 0;
        mem[604] <= 0;
        mem[605] <= 0;
        mem[606] <= 0;
        mem[607] <= 0;
        mem[608] <= 0;
        mem[609] <= 0;
        mem[610] <= 0;
        mem[611] <= 0;
        mem[612] <= 0;
        mem[613] <= 0;
        mem[614] <= 0;
        mem[615] <= 0;
        mem[616] <= 0;
        mem[617] <= 0;
        mem[618] <= 0;
        mem[619] <= 0;
        mem[620] <= 0;
        mem[621] <= 0;
        mem[622] <= 0;
        mem[623] <= 0;
        mem[624] <= 0;
        mem[625] <= 0;
        mem[626] <= 0;
        mem[627] <= 0;
        mem[628] <= 0;
        mem[629] <= 0;
        mem[630] <= 0;
        mem[631] <= 0;
        mem[632] <= 0;
        mem[633] <= 0;
        mem[634] <= 0;
        mem[635] <= 0;
        mem[636] <= 0;
        mem[637] <= 0;
        mem[638] <= 0;
        mem[639] <= 0;
        mem[640] <= 0;
        mem[641] <= 0;
        mem[642] <= 0;
        mem[643] <= 0;
        mem[644] <= 0;
        mem[645] <= 0;
        mem[646] <= 0;
        mem[647] <= 0;
        mem[648] <= 0;
        mem[649] <= 0;
        mem[650] <= 0;
        mem[651] <= 0;
        mem[652] <= 0;
        mem[653] <= 0;
        mem[654] <= 0;
        mem[655] <= 0;
        mem[656] <= 0;
        mem[657] <= 0;
        mem[658] <= 0;
        mem[659] <= 0;
        mem[660] <= 0;
        mem[661] <= 0;
        mem[662] <= 0;
        mem[663] <= 0;
        mem[664] <= 0;
        mem[665] <= 0;
        mem[666] <= 0;
        mem[667] <= 0;
        mem[668] <= 0;
        mem[669] <= 0;
        mem[670] <= 0;
        mem[671] <= 0;
        mem[672] <= 0;
        mem[673] <= 0;
        mem[674] <= 0;
        mem[675] <= 0;
        mem[676] <= 0;
        mem[677] <= 0;
        mem[678] <= 0;
        mem[679] <= 0;
        mem[680] <= 0;
        mem[681] <= 0;
        mem[682] <= 0;
        mem[683] <= 0;
        mem[684] <= 0;
        mem[685] <= 0;
        mem[686] <= 0;
        mem[687] <= 0;
        mem[688] <= 0;
        mem[689] <= 0;
        mem[690] <= 0;
        mem[691] <= 0;
        mem[692] <= 0;
        mem[693] <= 0;
        mem[694] <= 0;
        mem[695] <= 0;
        mem[696] <= 0;
        mem[697] <= 0;
        mem[698] <= 0;
        mem[699] <= 0;
        mem[700] <= 0;
        mem[701] <= 0;
        mem[702] <= 0;
        mem[703] <= 0;
        mem[704] <= 0;
        mem[705] <= 0;
        mem[706] <= 0;
        mem[707] <= 0;
        mem[708] <= 0;
        mem[709] <= 0;
        mem[710] <= 0;
        mem[711] <= 0;
        mem[712] <= 0;
        mem[713] <= 0;
        mem[714] <= 0;
        mem[715] <= 0;
        mem[716] <= 0;
        mem[717] <= 0;
        mem[718] <= 0;
        mem[719] <= 0;
        mem[720] <= 0;
        mem[721] <= 0;
        mem[722] <= 0;
        mem[723] <= 0;
        mem[724] <= 0;
        mem[725] <= 0;
        mem[726] <= 0;
        mem[727] <= 0;
        mem[728] <= 0;
        mem[729] <= 0;
        mem[730] <= 0;
        mem[731] <= 0;
        mem[732] <= 0;
        mem[733] <= 0;
        mem[734] <= 0;
        mem[735] <= 0;
        mem[736] <= 0;
        mem[737] <= 0;
        mem[738] <= 0;
        mem[739] <= 0;
        mem[740] <= 0;
        mem[741] <= 0;
        mem[742] <= 0;
        mem[743] <= 0;
        mem[744] <= 0;
        mem[745] <= 0;
        mem[746] <= 0;
        mem[747] <= 0;
        mem[748] <= 0;
        mem[749] <= 0;
        mem[750] <= 0;
        mem[751] <= 0;
        mem[752] <= 0;
        mem[753] <= 0;
        mem[754] <= 0;
        mem[755] <= 0;
        mem[756] <= 0;
        mem[757] <= 0;
        mem[758] <= 0;
        mem[759] <= 0;
        mem[760] <= 0;
        mem[761] <= 0;
        mem[762] <= 0;
        mem[763] <= 0;
        mem[764] <= 0;
        mem[765] <= 0;
        mem[766] <= 0;
        mem[767] <= 0;
        mem[768] <= 0;
        mem[769] <= 0;
        mem[770] <= 0;
        mem[771] <= 0;
        mem[772] <= 0;
        mem[773] <= 0;
        mem[774] <= 0;
        mem[775] <= 0;
        mem[776] <= 0;
        mem[777] <= 0;
        mem[778] <= 0;
        mem[779] <= 0;
        mem[780] <= 0;
        mem[781] <= 0;
        mem[782] <= 0;
        mem[783] <= 0;
        mem[784] <= 0;
        mem[785] <= 0;
        mem[786] <= 0;
        mem[787] <= 0;
        mem[788] <= 0;
        mem[789] <= 0;
        mem[790] <= 0;
        mem[791] <= 0;
        mem[792] <= 0;
        mem[793] <= 0;
        mem[794] <= 0;
        mem[795] <= 0;
        mem[796] <= 0;
        mem[797] <= 0;
        mem[798] <= 0;
        mem[799] <= 0;
        mem[800] <= 0;
        mem[801] <= 0;
        mem[802] <= 0;
        mem[803] <= 0;
        mem[804] <= 0;
        mem[805] <= 0;
        mem[806] <= 0;
        mem[807] <= 0;
        mem[808] <= 0;
        mem[809] <= 0;
        mem[810] <= 0;
        mem[811] <= 0;
        mem[812] <= 0;
        mem[813] <= 0;
        mem[814] <= 0;
        mem[815] <= 0;
        mem[816] <= 0;
        mem[817] <= 0;
        mem[818] <= 0;
        mem[819] <= 0;
        mem[820] <= 0;
        mem[821] <= 0;
        mem[822] <= 0;
        mem[823] <= 0;
        mem[824] <= 0;
        mem[825] <= 0;
        mem[826] <= 0;
        mem[827] <= 0;
        mem[828] <= 0;
        mem[829] <= 0;
        mem[830] <= 0;
        mem[831] <= 0;
        mem[832] <= 0;
        mem[833] <= 0;
        mem[834] <= 0;
        mem[835] <= 0;
        mem[836] <= 0;
        mem[837] <= 0;
        mem[838] <= 0;
        mem[839] <= 0;
        mem[840] <= 0;
        mem[841] <= 0;
        mem[842] <= 0;
        mem[843] <= 0;
        mem[844] <= 0;
        mem[845] <= 0;
        mem[846] <= 0;
        mem[847] <= 0;
        mem[848] <= 0;
        mem[849] <= 0;
        mem[850] <= 0;
        mem[851] <= 0;
        mem[852] <= 0;
        mem[853] <= 0;
        mem[854] <= 0;
        mem[855] <= 0;
        mem[856] <= 0;
        mem[857] <= 0;
        mem[858] <= 0;
        mem[859] <= 0;
        mem[860] <= 0;
        mem[861] <= 0;
        mem[862] <= 0;
        mem[863] <= 0;
        mem[864] <= 0;
        mem[865] <= 0;
        mem[866] <= 0;
        mem[867] <= 0;
        mem[868] <= 0;
        mem[869] <= 0;
        mem[870] <= 0;
        mem[871] <= 0;
        mem[872] <= 0;
        mem[873] <= 0;
        mem[874] <= 0;
        mem[875] <= 0;
        mem[876] <= 0;
        mem[877] <= 0;
        mem[878] <= 0;
        mem[879] <= 0;
        mem[880] <= 0;
        mem[881] <= 0;
        mem[882] <= 0;
        mem[883] <= 0;
        mem[884] <= 0;
        mem[885] <= 0;
        mem[886] <= 0;
        mem[887] <= 0;
        mem[888] <= 0;
        mem[889] <= 0;
        mem[890] <= 0;
        mem[891] <= 0;
        mem[892] <= 0;
        mem[893] <= 0;
        mem[894] <= 0;
        mem[895] <= 0;
        mem[896] <= 0;
        mem[897] <= 0;
        mem[898] <= 0;
        mem[899] <= 0;
        mem[900] <= 0;
        mem[901] <= 0;
        mem[902] <= 0;
        mem[903] <= 0;
        mem[904] <= 0;
        mem[905] <= 0;
        mem[906] <= 0;
        mem[907] <= 0;
        mem[908] <= 0;
        mem[909] <= 0;
        mem[910] <= 0;
        mem[911] <= 0;
        mem[912] <= 0;
        mem[913] <= 0;
        mem[914] <= 0;
        mem[915] <= 0;
        mem[916] <= 0;
        mem[917] <= 0;
        mem[918] <= 0;
        mem[919] <= 0;
        mem[920] <= 0;
        mem[921] <= 0;
        mem[922] <= 0;
        mem[923] <= 0;
        mem[924] <= 0;
        mem[925] <= 0;
        mem[926] <= 0;
        mem[927] <= 0;
        mem[928] <= 0;
        mem[929] <= 0;
        mem[930] <= 0;
        mem[931] <= 0;
        mem[932] <= 0;
        mem[933] <= 0;
        mem[934] <= 0;
        mem[935] <= 0;
        mem[936] <= 0;
        mem[937] <= 0;
        mem[938] <= 0;
        mem[939] <= 0;
        mem[940] <= 0;
        mem[941] <= 0;
        mem[942] <= 0;
        mem[943] <= 0;
        mem[944] <= 0;
        mem[945] <= 0;
        mem[946] <= 0;
        mem[947] <= 0;
        mem[948] <= 0;
        mem[949] <= 0;
        mem[950] <= 0;
        mem[951] <= 0;
        mem[952] <= 0;
        mem[953] <= 0;
        mem[954] <= 0;
        mem[955] <= 0;
        mem[956] <= 0;
        mem[957] <= 0;
        mem[958] <= 0;
        mem[959] <= 0;
        mem[960] <= 0;
        mem[961] <= 0;
        mem[962] <= 0;
        mem[963] <= 0;
        mem[964] <= 0;
        mem[965] <= 0;
        mem[966] <= 0;
        mem[967] <= 0;
        mem[968] <= 0;
        mem[969] <= 0;
        mem[970] <= 0;
        mem[971] <= 0;
        mem[972] <= 0;
        mem[973] <= 0;
        mem[974] <= 0;
        mem[975] <= 0;
        mem[976] <= 0;
        mem[977] <= 0;
        mem[978] <= 0;
        mem[979] <= 0;
        mem[980] <= 0;
        mem[981] <= 0;
        mem[982] <= 0;
        mem[983] <= 0;
        mem[984] <= 0;
        mem[985] <= 0;
        mem[986] <= 0;
        mem[987] <= 0;
        mem[988] <= 0;
        mem[989] <= 0;
        mem[990] <= 0;
        mem[991] <= 0;
        mem[992] <= 0;
        mem[993] <= 0;
        mem[994] <= 0;
        mem[995] <= 0;
        mem[996] <= 0;
        mem[997] <= 0;
        mem[998] <= 0;
        mem[999] <= 0;
        mem[1000] <= 0;
        mem[1001] <= 0;
        mem[1002] <= 0;
        mem[1003] <= 0;
        mem[1004] <= 0;
        mem[1005] <= 0;
        mem[1006] <= 0;
        mem[1007] <= 0;
        mem[1008] <= 0;
        mem[1009] <= 0;
        mem[1010] <= 0;
        mem[1011] <= 0;
        mem[1012] <= 0;
        mem[1013] <= 0;
        mem[1014] <= 0;
        mem[1015] <= 0;
        mem[1016] <= 0;
        mem[1017] <= 0;
        mem[1018] <= 0;
        mem[1019] <= 0;
        mem[1020] <= 0;
        mem[1021] <= 0;
        mem[1022] <= 0;
        mem[1023] <= 0;
    end
    else begin
        if ((i_mem_wr == 1)) begin
            if ((i_byte_wr == 1)) begin
                mem[i_address][8-1:0] <= i_wr_data[8-1:0];
            end
            else if ((i_2byte_wr == 1)) begin
                mem[i_address][16-1:0] <= i_wr_data[16-1:0];
            end
            else if ((i_4byte_wr == 1)) begin
                mem[i_address] <= i_wr_data;
            end
        end
    end
end


always @(i_se_mem_rd, i_mem_rd, i_4byte_rd, mem[0], mem[1], mem[2], mem[3], mem[4], mem[5], mem[6], mem[7], mem[8], mem[9], mem[10], mem[11], mem[12], mem[13], mem[14], mem[15], mem[16], mem[17], mem[18], mem[19], mem[20], mem[21], mem[22], mem[23], mem[24], mem[25], mem[26], mem[27], mem[28], mem[29], mem[30], mem[31], mem[32], mem[33], mem[34], mem[35], mem[36], mem[37], mem[38], mem[39], mem[40], mem[41], mem[42], mem[43], mem[44], mem[45], mem[46], mem[47], mem[48], mem[49], mem[50], mem[51], mem[52], mem[53], mem[54], mem[55], mem[56], mem[57], mem[58], mem[59], mem[60], mem[61], mem[62], mem[63], mem[64], mem[65], mem[66], mem[67], mem[68], mem[69], mem[70], mem[71], mem[72], mem[73], mem[74], mem[75], mem[76], mem[77], mem[78], mem[79], mem[80], mem[81], mem[82], mem[83], mem[84], mem[85], mem[86], mem[87], mem[88], mem[89], mem[90], mem[91], mem[92], mem[93], mem[94], mem[95], mem[96], mem[97], mem[98], mem[99], mem[100], mem[101], mem[102], mem[103], mem[104], mem[105], mem[106], mem[107], mem[108], mem[109], mem[110], mem[111], mem[112], mem[113], mem[114], mem[115], mem[116], mem[117], mem[118], mem[119], mem[120], mem[121], mem[122], mem[123], mem[124], mem[125], mem[126], mem[127], mem[128], mem[129], mem[130], mem[131], mem[132], mem[133], mem[134], mem[135], mem[136], mem[137], mem[138], mem[139], mem[140], mem[141], mem[142], mem[143], mem[144], mem[145], mem[146], mem[147], mem[148], mem[149], mem[150], mem[151], mem[152], mem[153], mem[154], mem[155], mem[156], mem[157], mem[158], mem[159], mem[160], mem[161], mem[162], mem[163], mem[164], mem[165], mem[166], mem[167], mem[168], mem[169], mem[170], mem[171], mem[172], mem[173], mem[174], mem[175], mem[176], mem[177], mem[178], mem[179], mem[180], mem[181], mem[182], mem[183], mem[184], mem[185], mem[186], mem[187], mem[188], mem[189], mem[190], mem[191], mem[192], mem[193], mem[194], mem[195], mem[196], mem[197], mem[198], mem[199], mem[200], mem[201], mem[202], mem[203], mem[204], mem[205], mem[206], mem[207], mem[208], mem[209], mem[210], mem[211], mem[212], mem[213], mem[214], mem[215], mem[216], mem[217], mem[218], mem[219], mem[220], mem[221], mem[222], mem[223], mem[224], mem[225], mem[226], mem[227], mem[228], mem[229], mem[230], mem[231], mem[232], mem[233], mem[234], mem[235], mem[236], mem[237], mem[238], mem[239], mem[240], mem[241], mem[242], mem[243], mem[244], mem[245], mem[246], mem[247], mem[248], mem[249], mem[250], mem[251], mem[252], mem[253], mem[254], mem[255], mem[256], mem[257], mem[258], mem[259], mem[260], mem[261], mem[262], mem[263], mem[264], mem[265], mem[266], mem[267], mem[268], mem[269], mem[270], mem[271], mem[272], mem[273], mem[274], mem[275], mem[276], mem[277], mem[278], mem[279], mem[280], mem[281], mem[282], mem[283], mem[284], mem[285], mem[286], mem[287], mem[288], mem[289], mem[290], mem[291], mem[292], mem[293], mem[294], mem[295], mem[296], mem[297], mem[298], mem[299], mem[300], mem[301], mem[302], mem[303], mem[304], mem[305], mem[306], mem[307], mem[308], mem[309], mem[310], mem[311], mem[312], mem[313], mem[314], mem[315], mem[316], mem[317], mem[318], mem[319], mem[320], mem[321], mem[322], mem[323], mem[324], mem[325], mem[326], mem[327], mem[328], mem[329], mem[330], mem[331], mem[332], mem[333], mem[334], mem[335], mem[336], mem[337], mem[338], mem[339], mem[340], mem[341], mem[342], mem[343], mem[344], mem[345], mem[346], mem[347], mem[348], mem[349], mem[350], mem[351], mem[352], mem[353], mem[354], mem[355], mem[356], mem[357], mem[358], mem[359], mem[360], mem[361], mem[362], mem[363], mem[364], mem[365], mem[366], mem[367], mem[368], mem[369], mem[370], mem[371], mem[372], mem[373], mem[374], mem[375], mem[376], mem[377], mem[378], mem[379], mem[380], mem[381], mem[382], mem[383], mem[384], mem[385], mem[386], mem[387], mem[388], mem[389], mem[390], mem[391], mem[392], mem[393], mem[394], mem[395], mem[396], mem[397], mem[398], mem[399], mem[400], mem[401], mem[402], mem[403], mem[404], mem[405], mem[406], mem[407], mem[408], mem[409], mem[410], mem[411], mem[412], mem[413], mem[414], mem[415], mem[416], mem[417], mem[418], mem[419], mem[420], mem[421], mem[422], mem[423], mem[424], mem[425], mem[426], mem[427], mem[428], mem[429], mem[430], mem[431], mem[432], mem[433], mem[434], mem[435], mem[436], mem[437], mem[438], mem[439], mem[440], mem[441], mem[442], mem[443], mem[444], mem[445], mem[446], mem[447], mem[448], mem[449], mem[450], mem[451], mem[452], mem[453], mem[454], mem[455], mem[456], mem[457], mem[458], mem[459], mem[460], mem[461], mem[462], mem[463], mem[464], mem[465], mem[466], mem[467], mem[468], mem[469], mem[470], mem[471], mem[472], mem[473], mem[474], mem[475], mem[476], mem[477], mem[478], mem[479], mem[480], mem[481], mem[482], mem[483], mem[484], mem[485], mem[486], mem[487], mem[488], mem[489], mem[490], mem[491], mem[492], mem[493], mem[494], mem[495], mem[496], mem[497], mem[498], mem[499], mem[500], mem[501], mem[502], mem[503], mem[504], mem[505], mem[506], mem[507], mem[508], mem[509], mem[510], mem[511], mem[512], mem[513], mem[514], mem[515], mem[516], mem[517], mem[518], mem[519], mem[520], mem[521], mem[522], mem[523], mem[524], mem[525], mem[526], mem[527], mem[528], mem[529], mem[530], mem[531], mem[532], mem[533], mem[534], mem[535], mem[536], mem[537], mem[538], mem[539], mem[540], mem[541], mem[542], mem[543], mem[544], mem[545], mem[546], mem[547], mem[548], mem[549], mem[550], mem[551], mem[552], mem[553], mem[554], mem[555], mem[556], mem[557], mem[558], mem[559], mem[560], mem[561], mem[562], mem[563], mem[564], mem[565], mem[566], mem[567], mem[568], mem[569], mem[570], mem[571], mem[572], mem[573], mem[574], mem[575], mem[576], mem[577], mem[578], mem[579], mem[580], mem[581], mem[582], mem[583], mem[584], mem[585], mem[586], mem[587], mem[588], mem[589], mem[590], mem[591], mem[592], mem[593], mem[594], mem[595], mem[596], mem[597], mem[598], mem[599], mem[600], mem[601], mem[602], mem[603], mem[604], mem[605], mem[606], mem[607], mem[608], mem[609], mem[610], mem[611], mem[612], mem[613], mem[614], mem[615], mem[616], mem[617], mem[618], mem[619], mem[620], mem[621], mem[622], mem[623], mem[624], mem[625], mem[626], mem[627], mem[628], mem[629], mem[630], mem[631], mem[632], mem[633], mem[634], mem[635], mem[636], mem[637], mem[638], mem[639], mem[640], mem[641], mem[642], mem[643], mem[644], mem[645], mem[646], mem[647], mem[648], mem[649], mem[650], mem[651], mem[652], mem[653], mem[654], mem[655], mem[656], mem[657], mem[658], mem[659], mem[660], mem[661], mem[662], mem[663], mem[664], mem[665], mem[666], mem[667], mem[668], mem[669], mem[670], mem[671], mem[672], mem[673], mem[674], mem[675], mem[676], mem[677], mem[678], mem[679], mem[680], mem[681], mem[682], mem[683], mem[684], mem[685], mem[686], mem[687], mem[688], mem[689], mem[690], mem[691], mem[692], mem[693], mem[694], mem[695], mem[696], mem[697], mem[698], mem[699], mem[700], mem[701], mem[702], mem[703], mem[704], mem[705], mem[706], mem[707], mem[708], mem[709], mem[710], mem[711], mem[712], mem[713], mem[714], mem[715], mem[716], mem[717], mem[718], mem[719], mem[720], mem[721], mem[722], mem[723], mem[724], mem[725], mem[726], mem[727], mem[728], mem[729], mem[730], mem[731], mem[732], mem[733], mem[734], mem[735], mem[736], mem[737], mem[738], mem[739], mem[740], mem[741], mem[742], mem[743], mem[744], mem[745], mem[746], mem[747], mem[748], mem[749], mem[750], mem[751], mem[752], mem[753], mem[754], mem[755], mem[756], mem[757], mem[758], mem[759], mem[760], mem[761], mem[762], mem[763], mem[764], mem[765], mem[766], mem[767], mem[768], mem[769], mem[770], mem[771], mem[772], mem[773], mem[774], mem[775], mem[776], mem[777], mem[778], mem[779], mem[780], mem[781], mem[782], mem[783], mem[784], mem[785], mem[786], mem[787], mem[788], mem[789], mem[790], mem[791], mem[792], mem[793], mem[794], mem[795], mem[796], mem[797], mem[798], mem[799], mem[800], mem[801], mem[802], mem[803], mem[804], mem[805], mem[806], mem[807], mem[808], mem[809], mem[810], mem[811], mem[812], mem[813], mem[814], mem[815], mem[816], mem[817], mem[818], mem[819], mem[820], mem[821], mem[822], mem[823], mem[824], mem[825], mem[826], mem[827], mem[828], mem[829], mem[830], mem[831], mem[832], mem[833], mem[834], mem[835], mem[836], mem[837], mem[838], mem[839], mem[840], mem[841], mem[842], mem[843], mem[844], mem[845], mem[846], mem[847], mem[848], mem[849], mem[850], mem[851], mem[852], mem[853], mem[854], mem[855], mem[856], mem[857], mem[858], mem[859], mem[860], mem[861], mem[862], mem[863], mem[864], mem[865], mem[866], mem[867], mem[868], mem[869], mem[870], mem[871], mem[872], mem[873], mem[874], mem[875], mem[876], mem[877], mem[878], mem[879], mem[880], mem[881], mem[882], mem[883], mem[884], mem[885], mem[886], mem[887], mem[888], mem[889], mem[890], mem[891], mem[892], mem[893], mem[894], mem[895], mem[896], mem[897], mem[898], mem[899], mem[900], mem[901], mem[902], mem[903], mem[904], mem[905], mem[906], mem[907], mem[908], mem[909], mem[910], mem[911], mem[912], mem[913], mem[914], mem[915], mem[916], mem[917], mem[918], mem[919], mem[920], mem[921], mem[922], mem[923], mem[924], mem[925], mem[926], mem[927], mem[928], mem[929], mem[930], mem[931], mem[932], mem[933], mem[934], mem[935], mem[936], mem[937], mem[938], mem[939], mem[940], mem[941], mem[942], mem[943], mem[944], mem[945], mem[946], mem[947], mem[948], mem[949], mem[950], mem[951], mem[952], mem[953], mem[954], mem[955], mem[956], mem[957], mem[958], mem[959], mem[960], mem[961], mem[962], mem[963], mem[964], mem[965], mem[966], mem[967], mem[968], mem[969], mem[970], mem[971], mem[972], mem[973], mem[974], mem[975], mem[976], mem[977], mem[978], mem[979], mem[980], mem[981], mem[982], mem[983], mem[984], mem[985], mem[986], mem[987], mem[988], mem[989], mem[990], mem[991], mem[992], mem[993], mem[994], mem[995], mem[996], mem[997], mem[998], mem[999], mem[1000], mem[1001], mem[1002], mem[1003], mem[1004], mem[1005], mem[1006], mem[1007], mem[1008], mem[1009], mem[1010], mem[1011], mem[1012], mem[1013], mem[1014], mem[1015], mem[1016], mem[1017], mem[1018], mem[1019], mem[1020], mem[1021], mem[1022], mem[1023], w_rd_data_2byte, i_address, w_rd_data_byte, i_byte_rd, i_2byte_rd) begin: DM_READ_LOGIC_1
    w_rd_data_byte = 0;
    w_rd_data_2byte = 0;
    w_rd_data = 0;
    if ((i_mem_rd == 1)) begin
        if ((i_byte_rd == 1)) begin
            w_rd_data_byte = mem[i_address][8-1:0];
            if ((i_se_mem_rd == 1)) begin
                w_rd_data = $signed(w_rd_data_byte);
            end
            else begin
                w_rd_data = {25'h0, w_rd_data_byte};
            end
        end
        else if ((i_2byte_rd == 1)) begin
            w_rd_data_2byte = mem[i_address][16-1:0];
            if ((i_se_mem_rd == 1)) begin
                w_rd_data = $signed(w_rd_data_2byte);
            end
            else begin
                w_rd_data = {17'h0, w_rd_data_2byte};
            end
        end
        else if ((i_4byte_rd == 1)) begin
            w_rd_data = mem[i_address];
        end
    end
end



assign o_rd_data = w_rd_data;

endmodule
